`ifndef MAC_TESTS_SVH
`define MAC_TESTS_SVH

`include "mac_base_test.sv"
`include "mac_small_packet_test.sv"
`include "mac_large_packet_test.sv"
`include "mac_oversized_packet_test.sv"
`include "mac_ipg_packet_test.sv"

`endif // MAC_TESTS_SVH

