`ifndef MAC_PKG_SV
`define MAC_PKG_SV
package mac_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "mac_transaction.sv"
  `include "mac_define.svh"
  `include "mac_driver.sv"
  `include "mac_monitor.sv"
  `include "mac_sequencer.sv"
  `include "mac_mst_driver.sv"
  `include "mac_mst_monitor.sv"
  `include "mac_mst_sequencer.sv"
  `include "mac_slv_monitor.sv"
  `include "mac_mst_agent.sv"
  `include "mac_slv_agent.sv"
endpackage


`endif
