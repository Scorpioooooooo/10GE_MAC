`ifndef MAC_SEQ_LIB_SVH
`define MAC_SEQ_LIB_SVH

`include "mac_base_element_sequence.sv"
`include "mac_reset_sequence.sv"
`include "mac_base_virtual_sequence.sv"
`include "mac_small_packet_virt_sequence.sv"
`include "mac_large_packet_virt_sequence.sv"
`include "mac_oversized_packet_virt_sequence.sv"
`include "mac_ipg_packet_virt_sequence.sv"


`endif
