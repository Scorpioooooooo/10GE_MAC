// pkt_tx_val
`define YES 1
`define NO 0

